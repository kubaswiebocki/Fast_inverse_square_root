`timescale 1ns / 1ps

//Ports and Register + Params
//////////////////////////////////////////////////////////////////////////////////
module TestBench_InvSqRoot;

reg clk;
reg rst = 0;
reg [31:0] DataIn;
wire [31:0] DataOut;

real DataOut_real;
reg [31:0] memory [0:99]; 
//////////////////////////////////////////////////////////////////////////////////

// Instantiate the InvertSQRoot module.
//////////////////////////////////////////////////////////////////////////////////
InvertSQRoot InvertSQRoot(
.DataOut(DataOut),

.clk(clk),
.rst(rst),
.DataIn(DataIn)
);
//////////////////////////////////////////////////////////////////////////////////

//Generate CLK
//////////////////////////////////////////////////////////////////////////////////
always begin
    clk = 1'b0;
    //DataOut_real =(2**(DataOut[30:23]-127))*($itor({1'b1,DataOut[22:0]})/2**23)*((-1)**(DataOut[31]));
    #5;
    clk = 1'b1;
    #5; 
    end
    
//////////////////////////////////////////////////////////////////////////////////

//Command window
//////////////////////////////////////////////////////////////////////////////////
integer i;

initial begin
    $readmemb("InputData.mem", memory);
    for (i=0; i<100; i=i+1) begin
        DataIn = memory[i];
        #10;
        end
    $display("Simulation is over, check the waveforms.");
    $stop;
    end
//////////////////////////////////////////////////////////////////////////////////

endmodule