`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Lukasz Orzel
// Engineer: Jakub Swiebocki
// Module Name: InvertSQRoot
// Project Name: Fast inverse square root 
// Target Devices: ZedBoard
// Tool Versions: Vivado 2018.2
// 
//////////////////////////////////////////////////////////////////////////////////

//Conncet and Register + Params
//////////////////////////////////////////////////////////////////////////////////
module InvertSQRoot(
    output reg  [31:0] DataOut,
    
    input wire [31:0] DataIn,
    input wire clk,
    input wire rst
    );
    
reg  [31:0] Data_temp, Data_temp_nxt;
reg  [31:0] DataOut_nxt;
reg  [31:0] i, exponent;

localparam  E = 127;
localparam  MAGIC = 32'h5f3759df;

//////////////////////////////////////////////////////////////////////////////////

//Zegar
//////////////////////////////////////////////////////////////////////////////////
always@ (posedge clk) begin
    if(rst) begin
        DataOut <= 0;
        end
    else begin
        DataOut <= DataOut_nxt;
        Data_temp <= Data_temp_nxt;
        end
    end
//////////////////////////////////////////////////////////////////////////////////

//Algorytm InverSQRoot
//////////////////////////////////////////////////////////////////////////////////
always@* begin
    DataOut_nxt = MAGIC - (DataIn >> 1);    
end
//////////////////////////////////////////////////////////////////////////////////
endmodule
