`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Łukasz Orzeł
// Engineer: Jakub Świebocki
// Module Name: InvertSQRoot
// Project Name: Fast inverse square root 
// Target Devices: ZedBoard
// Tool Versions: Vivado 2018.2
// 
//////////////////////////////////////////////////////////////////////////////////


module InvertSQRoot(

    );
endmodule
