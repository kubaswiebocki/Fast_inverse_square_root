`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Lukasz Orzel�
// Engineer: Jakub Swiebocki
// Module Name: InvertSQRoot
// Project Name: Fast inverse square root 
// Target Devices: ZedBoard
// Tool Versions: Vivado 2018.2
// 
//////////////////////////////////////////////////////////////////////////////////

//Conncet and Register + Params
//////////////////////////////////////////////////////////////////////////////////
module InvertSQRoot(
    output reg  [31:0] DataOut,
    
    input wire [31:0] DataIn,
    input wire clk,
    input wire rst
    );
    
reg  [31:0] Data_temp, Data_temp_nxt;
reg  [31:0] DataOut_nxt;

localparam FXPratio = 1024;
//////////////////////////////////////////////////////////////////////////////////

//Zegar
//////////////////////////////////////////////////////////////////////////////////
always@ (posedge clk) begin
    if(rst) begin
        DataOut <= 0;
        end
    else begin
        DataOut <= DataOut_nxt;
        Data_temp <= Data_temp_nxt;
        end
    end
//////////////////////////////////////////////////////////////////////////////////

//Algorytm InverSQRoot
//////////////////////////////////////////////////////////////////////////////////
always@* begin
    Data_temp_nxt <= DataIn*FXPratio ;
    DataOut_nxt <= 32'h5F3759DF - (DataIn>>1);
    end
//////////////////////////////////////////////////////////////////////////////////

endmodule
